class MyTransaction extends  uvm_sequence_item;
	

endclass